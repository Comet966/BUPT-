﻿//四位串行加法器module key_1 (    input clk,       input [3:0] key,    input [3:0] sw,        output [8:0] seg1,	 output [8:0] seg2,	 output [7:0] led);wire key1_on;wire key2_on;wire key3_on;wire [3:0] sum_wire;wire cout_wire;reg [1:0] state;reg [3:0] num1;reg [3:0] num2;reg [7:0] num3;reg [8:0] seg1_value;reg [8:0] seg2_value;reg [3:0] sw_value;reg [7:0] led_value;reg cin;initial beginstate = 2'b00;num1 = 4'b0000;num2 = 4'b0000;led_value = ~8'b1111_1111;cin = 1'b0;endassign led = ~led_value;assign seg2 = seg1_value;assign seg1 = seg2_value;serial_adder_4bit add_4bit(.a(num1),.b(num2),.cin(cin),.sum(sum_wire),.cout(cout_wire));always @(posedge clk)beginsw_value <= {sw[0], sw[1], sw[2], sw[3]};if(key[0] == 0)beginnum1 <= sw_value;state <= 2'b01;led_value[0] <= state[0];led_value[1] <= state[1];//0~15译码器case(num1)4'h0:begin seg1_value<=9'h3f;seg2_value<=9'h3f;end4'h1:begin seg1_value<=9'h06;seg2_value<=9'h3f;end 4'h2:begin seg1_value<=9'h5b;seg2_value<=9'h3f;end4'h3:begin seg1_value<=9'h4f;seg2_value<=9'h3f;end4'h4:begin seg1_value<=9'h66;seg2_value<=9'h3f;end   4'h5:begin seg1_value<=9'h6d;seg2_value<=9'h3f;end  4'h6:begin seg1_value<=9'h7d;seg2_value<=9'h3f;end4'h7:begin seg1_value<=9'h07;seg2_value<=9'h3f;end4'h8:begin seg1_value<=9'h7f;seg2_value<=9'h3f;end4'h9:begin seg1_value<=9'h6f;seg2_value<=9'h3f;end4'hA:begin seg1_value<=9'h3f;seg2_value<=9'h06;end4'hB:begin seg1_value<=9'h06;seg2_value<=9'h06;end 4'hC:begin seg1_value<=9'h5b;seg2_value<=9'h06;end4'hD:begin seg1_value<=9'h4f;seg2_value<=9'h06;end4'hE:begin seg1_value<=9'h66;seg2_value<=9'h06;end   4'hF:begin seg1_value<=9'h6d;seg2_value<=9'h06;end  default:begin  seg1_value<=9'h3f;seg2_value<=9'h3f;endendcaseendif(key[1] == 0)beginnum2 <= sw_value;state <= 2'b11;led_value[0] <= state[0];led_value[1] <= state[1];case(num2)4'h0:begin seg1_value<=9'h3f;seg2_value<=9'h3f;end4'h1:begin seg1_value<=9'h06;seg2_value<=9'h3f;end 4'h2:begin seg1_value<=9'h5b;seg2_value<=9'h3f;end4'h3:begin seg1_value<=9'h4f;seg2_value<=9'h3f;end4'h4:begin seg1_value<=9'h66;seg2_value<=9'h3f;end   4'h5:begin seg1_value<=9'h6d;seg2_value<=9'h3f;end  4'h6:begin seg1_value<=9'h7d;seg2_value<=9'h3f;end4'h7:begin seg1_value<=9'h07;seg2_value<=9'h3f;end4'h8:begin seg1_value<=9'h7f;seg2_value<=9'h3f;end4'h9:begin seg1_value<=9'h6f;seg2_value<=9'h3f;end4'hA:begin seg1_value<=9'h3f;seg2_value<=9'h06;end4'hB:begin seg1_value<=9'h06;seg2_value<=9'h06;end 4'hC:begin seg1_value<=9'h5b;seg2_value<=9'h06;end4'hD:begin seg1_value<=9'h4f;seg2_value<=9'h06;end4'hE:begin seg1_value<=9'h66;seg2_value<=9'h06;end   4'hF:begin seg1_value<=9'h6d;seg2_value<=9'h06;end  default:begin  seg1_value<=9'h3f;seg2_value<=9'h3f;endendcaseendif(key[2] == 0)begin// num3 <= num1 + num2;num3 <= {cout_wire,sum_wire};state <= 2'b00;led_value[0] <= state[0];led_value[1] <= state[1];case(num3 % 4'hA)5'h0:seg1_value<=9'h3f;5'h1:seg1_value<=9'h06; 5'h2:seg1_value<=9'h5b;5'h3:seg1_value<=9'h4f;5'h4:seg1_value<=9'h66;   5'h5:seg1_value<=9'h6d;  5'h6:seg1_value<=9'h7d;5'h7:seg1_value<=9'h07;5'h8:seg1_value<=9'h7f;5'h9:seg1_value<=9'h6f;default: seg1_value<=9'h00;endcaseif(num3 < 5'd10)seg2_value<=9'h3f;else if(num3 <5'd20)seg2_value<=9'h06;else if(num3 < 5'd30)seg2_value<=9'h5b;else seg2_value<=9'h4f;endendendmodule