﻿module JK_trigger(J,K,clk,Q,Qn);
input J,K,clk;
output reg Q;
output wire Qn;
assign Qn = ~Q;
always@(posedge clk)
case({J,K})
2'b00:Q<=Q;
2'b01:Q<=1'b0;
2'b10:Q<=1'b1;
2'b11:Q<=~Q;
endcase

endmodule

module fpga_prj(clk,clr,oe,dout);
input wire clk,clr,oe;
output wire [3:0] dout;

wire [1:0]jk0,jk1,jk2,jk3;
wire q0,q1,q2,q3;

JK_trigger
jk0_inst(.J(1),.K(1),.clk(clk),.Q(q0),.Qn());
JK_trigger
jk1_inst(.J(q0),.K(1),.clk(clk),.Q(q1),.Qn());
JK_trigger
jk2_inst(.J(q1),.K(1),.clk(clk),.Q(q2),.Qn());
JK_trigger
jk3_inst(.J(q2),.K(1),.clk(clk),.Q(q3),.Qn());

assign jk0 = {q3,q2};
assign jk1 = {q3,q2};
assign jk2 = {q3,q2};
assign jk3 = {q3,q2};

assign dout = {q3,q2,q1,q0};
endmodule

