﻿//例化D触发器实现74HC595（四位并行移位寄存器）
module D_ff(D_in , clk , q , q_bar );
input D_in,clk;
output q,q_bar;
reg q_value;

always@(posedge clk)begin

q_value <= D_in;

end
endmodule

module fpga_prj(clk,x_in,q1,q2,q3,q4);
input clk,x_in;
output q1,q2,q3,q4;
D_ff D_ff1(.D_in(x_in),.clk(clk),.q(q1));
D_ff D_ff2(.D_in(q1),.clk(clk),.q(q2));
D_ff D_ff3(.D_in(q2),.clk(clk),.q(q3));
D_ff D_ff4(.D_in(q3),.clk(clk),.q(q4));

endmodule
