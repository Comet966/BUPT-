﻿module fadd(a, b, Cin, Cout, Sum);    input a, b, Cin;    output Sum, Cout;    assign {Cout, Sum} = a + b + Cin;endmodulemodule serial_adder_4bit(    input [3:0] a, b,  // 两组 4 位加数    input cin,         // 低位来的进位    output [3:0] sum,  // 加法运算的结果    output cout        // 最高位的进位);    wire [3:0] c;  // 进位线    fadd fa0(.a(a[0]), .b(b[0]), .Cin(cin),  .Sum(sum[0]), .Cout(c[0]));    fadd fa1(.a(a[1]), .b(b[1]), .Cin(c[0]), .Sum(sum[1]), .Cout(c[1]));    fadd fa2(.a(a[2]), .b(b[2]), .Cin(c[1]), .Sum(sum[2]), .Cout(c[2]));    fadd fa3(.a(a[3]), .b(b[3]), .Cin(c[2]), .Sum(sum[3]), .Cout(cout));endmodule