﻿//汽车尾灯控制module fpga_prj(clk,sw,rgb_1,rgb_2,seg1);input clk;input [2:0] sw;output rgb_1;output rgb_2;output [8:0] seg1;rgb(.clk(clk),.sig(sw),.out_rgb({rgb_1,rgb_2}));seg(.clk(clk),.seg(seg1),.sw({1'b0,sw}));endmodule//rgb闪烁模块sig为一位控制信号module rgb(clk,sig,out_rgb);input clk;input [2:0] sig;output [1:0] out_rgb;reg [1:0] rgb;reg [26:0] num;assign out_rgb = rgb;parameter count = 12_000_000;always@(posedge clk)beginnum<= num+1;if(num >= 12_000_000)begincase(sig)3'b001:rgb <= ~rgb;3'b010:rgb <= {~rgb[1],1'b1};3'b011:rgb <= {1'b1,~rgb[0]};3'b100:rgb <= 2'b00;default: rgb <= 2'b11;endcasenum <= 0;endendendmodulemodule seg(clk,seg,sw);input clk;input [3:0]sw;output [8:0]seg;reg [8:0] seg_value;assign seg = seg_value;always@(posedge clk)begincase(sw)4'h0:seg_value<=9'h3f;4'h1:seg_value<=9'h06; 4'h2:seg_value<=9'h5b;4'h3:seg_value<=9'h4f;4'h4:seg_value<=9'h66;   4'h5:seg_value<=9'h6d;  4'h6:seg_value<=9'h7d;4'h7:seg_value<=9'h07;4'h8:seg_value<=9'h7f;4'h9:seg_value<=9'h6f;default:seg_value <= seg_value;endcaseendendmodule