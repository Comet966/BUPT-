﻿module fpga_prj(    input wire clk,      // 时钟信号    input wire rst,      // 异步复位信号（高电平有效）    input wire data,     // 串行输入数据（1位）    output reg detected  // 输出信号：检测到"101"时为1);// 状态定义（使用参数，便于修改）parameter S0 = 2'b00;  // 初始状态parameter S1 = 2'b01;  // 检测到"1"parameter S2 = 2'b10;  // 检测到"10"parameter S3 = 2'b11;  // 检测到"101"// 状态寄存器（当前状态）reg [1:0] current_state, next_state;// 状态转移：时序逻辑（同步更新当前状态）always @(posedge clk or posedge rst) begin    if (rst) begin        current_state <= S0;  // 复位到初始状态    end else begin        current_state <= next_state;  // 更新状态    endend// 下一状态逻辑：组合逻辑always @(*) begin    case (current_state)        S0: begin            if (data == 1'b1) next_state = S1;            else next_state = S0;        end        S1: begin            if (data == 1'b0) next_state = S2;            else next_state = S1;        end        S2: begin            if (data == 1'b1) next_state = S3;            else next_state = S0;        end        S3: begin            next_state = S0;  // 序列检测后返回初始        end        default: next_state = S0;    endcaseend// 输出逻辑：Moore机（输出仅依赖当前状态）always @(*) begin    if (current_state == S3) detected = 1'b1;    else detected = 1'b0;endendmodule