﻿//使用例化译码器模块的方式实现BCD控制数码管

module fpga_prj(seg1,sw);
input [3:0] sw;
output [8:0] seg1;

seg_encoder en0(.num({sw[0],sw[1],sw[2],sw[3]}),.output_value(seg1));


endmodule



module seg_encoder(num,output_value);

input [3:0] num;
output reg [8:0] output_value;
always@(*)begin
case(num)
4'h0:output_value=9'h3f;
4'h1:output_value=9'h06; 
4'h2:output_value=9'h5b;
4'h3:output_value=9'h4f;
4'h4:output_value=9'h66;   
4'h5:output_value=9'h6d;  
4'h6:output_value=9'h7d;
4'h7:output_value=9'h07;
4'h8:output_value=9'h7f;
4'h9:output_value=9'h6f;
default: output_value=9'h00;

endcase
end
endmodule

